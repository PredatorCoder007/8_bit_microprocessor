//8-bit microprocessor design using VHDL

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity processor is
     
     Port ( clk : in STD_LOGIC;
            value : out STD_LOGIC_VECTOR(7 downto 0));

end processor

architecture Behavioral of processor is

begin

end Behavioral;